`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:06:35 01/19/2017 
// Design Name: 
// Module Name:    R4BoothMultiplier 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module R4BoothMultiplier(
    input [15:0] multiplicand,
    input [15:0] multiplier,
    output [31:0] product
    );


endmodule
